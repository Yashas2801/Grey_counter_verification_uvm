package grey_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "grey_xtn.sv"

  `include "grey_seqs.sv"

  `include "grey_driver.sv"
  `include "grey_moniter.sv"
  `include "grey_sequencer.sv"
  `include "grey_agent.sv"

  `include "grey_coverage.sv"
  `include "grey_env.sv"

  `include "grey_test.sv"
endpackage
